library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity cache_tb is 
end entity;

architecture behavioral of cache_tb is
    begin
    end architecture;