library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity exception is 
end entity;

architecture behavioral of exception is
    begin
    end architecture;