library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity gpio_peripheral is 
end entity;

architecture behavioral of gpio_peripheral is
    begin
    end architecture;