library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity reg is 
end entity;

architecture behavioral of reg is
    begin
    end architecture;