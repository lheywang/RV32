/*
 *  File :      rtl/rv32.sv
 *
 *  Author :    l.heywang <leonard.heywang@proton.me>
 *  Date :      
 *  
 *  Brief :     This file is the top level of the whole core.
 *              Feel free to modify it to get the right core for your needs !
 */

`timescale 1ns / 1ps

module rv32 ();

endmodule
;
