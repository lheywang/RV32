library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity rv32 is 
end entity;

architecture behavioral of rv32 is
    begin
    end architecture;