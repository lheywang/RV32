library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity exception_tb is 
end entity;

architecture behavioral of exception_tb is
    begin
    end architecture;