library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity memcontroller is 
end entity;

architecture behavioral of memcontroller is
    begin
    end architecture;