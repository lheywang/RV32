library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity sdram is 
end entity;

architecture behavioral of sdram is
    begin
    end architecture;