library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity i_decoder is 
end entity;

architecture behavioral of i_decoder is
    begin
    end architecture;