LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;

ENTITY gpio_peripheral IS
END ENTITY;

ARCHITECTURE behavioral OF gpio_peripheral IS
BEGIN
END ARCHITECTURE;