library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity memcontroller_tb is 
end entity;

architecture behavioral of memcontroller_tb is
    begin
    end architecture;