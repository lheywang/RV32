/*
 *  File :      rtl/core/assembly/assembly_csr.sv
 *
 *  Author :    l.heywang <leonard.heywang@proton.me>
 *  Date :      25/10.2025
 *  
 *  Brief :     This file assemble all of the CSR with it's associated
 *              counters. This make the global core assembly much
 *              more readable.
 */

module assembly_csr ();

endmodule
