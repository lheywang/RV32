library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity alu_tb is 
end entity;

architecture behavioral of alu_tb is
    begin
    end architecture;