library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.common.all;

entity decoder is 
    generic (
        XLEN :      integer := 32                                           -- Width of the data outputs. 
                                                                            -- Warning : This does not change the number of registers not i_instruction lenght
    );
    port (
        -- instruction input
        instruction :   in      std_logic_vector(31 downto 0);

        -- shift enable
        shift_en :      in      std_logic;

        -- outputs
        -- buses
        rs1 :           out     std_logic_vector((XLEN / 8) downto 0)                   := (others => '0');
        rs2 :           out     std_logic_vector((XLEN / 8) downto 0)                   := (others => '0');   
        rd :            out     std_logic_vector((XLEN / 8) downto 0)                   := (others => '0');
        imm :           out     std_logic_vector((XLEN - 1) downto 0)                   := (others => '0');
        opcode :        out     instructions;                         
        -- signals
        illegal :       out     std_logic;

        -- Clocks
        clock :         in      std_logic;
        clock_en :      in      std_logic;
        nRST :          in      std_logic
    );
end entity;

architecture behavioral of decoder is

        -- Defining the different selected_decoders
        type decocders_type is (U, I, R, B, S, J, default_t, illegal_t, NOP);

        -- signals
        signal illegal_internal :      std_logic                                        := '0';
        signal illegal_internal2 :     std_logic                                        := '0';
        signal illegal_internal_out :  std_logic                                        := '0';

        -- Internal states
        signal selected_decoder :      decocders_type                                   := default_t;

        -- Latchs outputs
        signal  rs1_internal :          std_logic_vector(4 downto 0)                    := (others => '0');
        signal  rs2_internal :          std_logic_vector(4 downto 0)                    := (others => '0');
        signal  rd_internal :           std_logic_vector(4 downto 0)                    := (others => '0');
        signal  imm_internal :          std_logic_vector((XLEN - 1) downto 0)           := (others => '0');

        -- Internal instruction bus, with the right endianess
        signal  i_instruction :         std_logic_vector(31 downto 0)                   := (others => '0');
        signal  r_instruction :         std_logic_vector(31 downto 0)                   := (others => '0');

        -- remove the first decoder cycle glitch
        signal  first_flag :            std_logic                                       := '0';

    begin

        -- Register the input, to enable constant delays between decoders outputs
        P0 : process(clock, nRST)
        begin
            if (nRST = '0') then
                r_instruction <= (others => '0');
                first_flag <= '0';

            elsif rising_edge(clock) and (clock_en = '1') and (shift_en = '1') then
                if (first_flag = '1') then
                    r_instruction <= instruction;
                else
                    first_flag <= '1';
                end if;

            end if;

        end process;

        -- Endianess correctors
        U1 : entity work.endianess(rtl)
            generic map (
                XLEN        =>  32
            )
            port map (
                datain      =>  r_instruction,
                dataout     =>  i_instruction
            );

        -- Combinantional decoder, select the wanted decoder
        -- Using this not synced to clock enable to split the logic in half, and reduce the critical path
        -- Before, we've got Fmax = ~100 MHz because of it's too long logic.
        -- After, quartus report Fmax = ~230 MHz, because of the middle registering process.
        P1 : process(nRST, i_instruction) 
            begin

                if (nRST = '0') then
                    illegal_internal    <= '0';
                    selected_decoder    <= default_t;

                else

                    -- Select the opcode, and perform an instruction size check (last two bits must be "11").
                    case i_instruction(6 downto 0) is

                        when "0110111" =>               -- LUI
                            selected_decoder <= U;
                            illegal_internal <= '0';
                        when "0010111" =>               -- AUIPC
                            selected_decoder <= U;
                            illegal_internal <= '0';

                        when "0010011" =>               -- Immediates
                            selected_decoder <= I;
                            illegal_internal <= '0';
                        when "0001111" =>               -- FENCE
                            selected_decoder <= I;
                            illegal_internal <= '0';
                        when "1100111" =>               --(JALR)
                            selected_decoder <= I;
                            illegal_internal <= '0';
                        when "1110011" =>               -- Calls
                            selected_decoder <= I;
                            illegal_internal <= '0';
                        when "0000011" =>               -- Store
                            selected_decoder <= I;
                            illegal_internal <= '0';

                        when "0110011" =>               -- Register operations
                            selected_decoder <= R;
                            illegal_internal <= '0';
                        
                        when "1100011" =>               -- Branchs
                            selected_decoder <= B;
                            illegal_internal <= '0';
                        
                        when "0100011" =>               -- Loads
                            selected_decoder <= S;
                            illegal_internal <= '0';

                        when "1101111" =>               -- Jumps
                            selected_decoder <= J;
                            illegal_internal <= '0';

                        when "0000000" =>               -- All zero, seen as NOP
                            selected_decoder <= NOP;
                            illegal_internal <= '0';

                        when others =>
                            selected_decoder <= illegal_t;
                            illegal_internal <= '1';

                    end case;
                end if;
                
            end process;

        -- P2 : process(clock, nRST, clock_en)
        --     begin
        --         if (nRST = '0') then    
        --             r_selected_decoder <= default_t;

        --         elsif rising_edge(clock) and (clock_en = '1') then
        --             r_selected_decoder <= selected_decoder;

        --         end if;
        --     end process;

        -- Hardware selected_decoder selection logic
        -- This process is actually clocked, because we need synchronous outputs.
        P3 : process(clock, clock_en, nRST)
            begin
                if (nRST = '0') then
                    rs1_internal <= (others => '0');
                    rs2_internal <= (others => '0');
                    imm_internal <= (others => '0');
                    rd_internal <= (others => '0');
                    opcode <= i_NOP;
                    illegal_internal2 <= '0';

                elsif rising_edge(clock) and (clock_en = '1') and (shift_en = '1') then

                    case selected_decoder is 

                        -- Register to register operation
                        when R =>
                            rd_internal <=                                  i_instruction(11 downto 7);
                            rs1_internal <=                                 i_instruction(19 downto 15);
                                                                           
                            rs2_internal <=                                 i_instruction(24 downto 20);
                            imm_internal <=                                 (others => '0');
                        
                            -- i_instruction identification
                            case i_instruction(31 downto 25) is 

                                when "0000000" => -- ADD SLL SLT XOR SRL OR AND

                                    case i_instruction(14 downto 12) is

                                        when "000" =>
                                            opcode <= i_ADD;
                                            illegal_internal2 <= '0';
                                        when "001" =>
                                            opcode <= i_SLL;
                                            illegal_internal2 <= '0';
                                        when "010" =>
                                            opcode <= i_SLT;
                                            illegal_internal2 <= '0';
                                        when "011" =>
                                            opcode <= i_SLTU;
                                            illegal_internal2 <= '0';
                                        when "100" =>
                                            opcode <= i_XOR;
                                            illegal_internal2 <= '0';
                                        when "101" =>
                                            opcode <= i_SRL;
                                            illegal_internal2 <= '0';
                                        when "110" => 
                                            opcode <= i_OR;
                                            illegal_internal2 <= '0';
                                        when "111" =>
                                            opcode <= i_AND; 
                                            illegal_internal2 <= '0';
                                        when others =>
                                            opcode <= i_NOP;
                                            illegal_internal2 <= '1';

                                    end case;

                                when "0100000" => -- SUB SRA

                                    case i_instruction(14 downto 12) is

                                        when "000" =>
                                            opcode <= i_SUB;
                                            illegal_internal2 <= '0';
                                        when "101" =>
                                            opcode <= i_SRA;
                                            illegal_internal2 <= '0';
                                        when others =>
                                            opcode <= i_NOP;
                                            illegal_internal2 <= '1';

                                    end case;

                                when others => 
                                    opcode <= i_NOP;
                                    illegal_internal2 <= '1';

                            end case;

                        -- Immediate to register operation
                        when I =>
                            rd_internal <=                                  i_instruction(11 downto 7);
                            rs1_internal <=                                 i_instruction(19 downto 15); 
                            rs2_internal <=                                 (others => '0');
                            imm_internal <=                                 (others => i_instruction(31));
                            imm_internal(11 downto 0) <=                    i_instruction(31 downto 20);
                            
                            -- i_instruction identification
                            case i_instruction(6 downto 2) is

                                when "00100" => 
                            
                                    case i_instruction(14 downto 12) is

                                        when "000" =>
                                            opcode <= i_ADDI;
                                            illegal_internal2 <= '0';
                                        when "001" =>
                                            opcode <= i_SLLI;
                                            illegal_internal2 <= '0';
                                        when "010" =>
                                            opcode <= i_SLTI;
                                            illegal_internal2 <= '0';
                                        when "011" =>
                                            opcode <= i_SLTIU;
                                            illegal_internal2 <= '0';
                                        when "100" =>
                                            opcode <= i_XORI;
                                            illegal_internal2 <= '0';
                                        when "110" =>
                                            opcode <= i_ORI;
                                            illegal_internal2 <= '0';
                                        when "101" => 
                                            if (i_instruction(30) = '1') then
                                                opcode <= i_SRAI;
                                                illegal_internal2 <= '0';
                                            else
                                                opcode <= i_SRLI;
                                                illegal_internal2 <= '0';
                                            end if;

                                        when "111" =>
                                            opcode <= i_ANDI; 
                                            illegal_internal2 <= '0';
                                        when others =>
                                            opcode <= i_NOP;
                                            illegal_internal2 <= '0';

                                    end case;
                                
                                when "00011" =>
                                    opcode <= i_FENCE; 
                                    illegal_internal2 <= '0';

                                when "00000" =>

                                    case i_instruction(14 downto 12) is

                                        when "000" =>
                                            opcode <= i_LB;
                                            illegal_internal2 <= '0';
                                        when "001" =>
                                            opcode <= i_LH;
                                            illegal_internal2 <= '0';
                                        when "010" =>
                                            opcode <= i_LW;
                                            illegal_internal2 <= '0';
                                        when "100" =>
                                            opcode <= i_LBU;
                                            illegal_internal2 <= '0';
                                        when "101" =>
                                            opcode <= i_LHU;
                                            illegal_internal2 <= '0';
                                        when others =>
                                            opcode <= i_NOP; 
                                            illegal_internal2 <= '1';

                                    end case;
                                        
                                when "11001" => 
                                    if (i_instruction(14 downto 12) = "000") then
                                        opcode <= i_JALR; 
                                        illegal_internal2 <= '0';
                                    else
                                        opcode <= i_NOP;
                                        illegal_internal2 <= '1';
                                    end if;

                                when "11100" =>

                                    case i_instruction(14 downto 12) is

                                        when "001" =>
                                            opcode <= i_CSRRW;
                                            illegal_internal2 <= '0';
                                        when "010" =>
                                            opcode <= i_CSRRS;
                                            illegal_internal2 <= '0';
                                        when "011" =>
                                            opcode <= i_CSRRC;
                                            illegal_internal2 <= '0';
                                        when "101" =>
                                            opcode <= i_CSRRWI;
                                            illegal_internal2 <= '0';
                                        when "110" =>
                                            opcode <= i_CSRRSI;
                                            illegal_internal2 <= '0';
                                        when "111" =>
                                            opcode <= i_CSRRCI;
                                            illegal_internal2 <= '0';
                                        when "000" =>

                                            case i_instruction(31 downto 20) is

                                                when X"000" =>
                                                    opcode <= i_ECALL;
                                                    illegal_internal2 <= '0';
                                                when X"001" =>
                                                    opcode <= i_EBREAK;
                                                    illegal_internal2 <= '0';
                                                when X"302" =>
                                                    opcode <= i_MRET;
                                                    illegal_internal2 <= '0';
                                                when others =>
                                                    opcode <= i_NOP;
                                                    illegal_internal2 <= '1';

                                            end case;

                                        when others =>
                                            opcode <= i_NOP; 
                                            illegal_internal2 <= '1';

                                    end case;

                                when others => 
                                    opcode <= i_NOP;
                                    illegal_internal2 <= '1';

                            end case;


                        -- Memory operation
                        when S =>
                            rd_internal <=                                  (others => '0');
                            rs1_internal <=                                 i_instruction(19 downto 15); 
                            rs2_internal <=                                 i_instruction(24 downto 20);
                            imm_internal <=                                 (others => i_instruction(31));
                            imm_internal(11 downto 0) <=                    i_instruction(31 downto 25)                       
                                                                          & i_instruction(11 downto 7);

                            -- i_instruction identification
                            case i_instruction(14 downto 12) is

                                when "000" =>
                                    opcode <= i_SB; 
                                    illegal_internal2 <= '0';
                                when "001" =>
                                    opcode <= i_SH; 
                                    illegal_internal2 <= '0';
                                when "010" =>
                                    opcode <= i_SW; 
                                    illegal_internal2 <= '0';
                                when others =>

                            end case;

                        -- Branches
                        when B =>
                            rd_internal <=                                  (others => '0');
                            rs1_internal <=                                 i_instruction(19 downto 15);
                            rs2_internal <=                                 i_instruction(24 downto 20);
                            imm_internal <=                                 (others => i_instruction(31));
                            imm_internal(11 downto 0) <=                    i_instruction(31)                                 
                                                                          & i_instruction(7)                
                                                                          & i_instruction(30 downto 25)         
                                                                          & i_instruction(11 downto 8);

                            -- i_instruction identification
                            case i_instruction(14 downto 12) is

                                when "000" =>
                                    opcode <= i_BEQ; 
                                    illegal_internal2 <= '0';
                                when "001" =>
                                    opcode <= i_BNE; 
                                    illegal_internal2 <= '0';
                                when "100" =>
                                    opcode <= i_BLT; 
                                    illegal_internal2 <= '0';
                                when "101" =>
                                    opcode <= i_BGE; 
                                    illegal_internal2 <= '0';
                                when "110" =>
                                    opcode <= i_BLTU; 
                                    illegal_internal2 <= '0';
                                when "111" =>
                                    opcode <= i_BGEU; 
                                    illegal_internal2 <= '0';
                                when others =>
                                    opcode <= i_NOP; 
                                    illegal_internal2 <= '1';

                            end case;

                        -- Immediates values loading
                        when U =>
                            rd_internal <=                                   i_instruction(11 downto 7);
                            rs1_internal <=                                  (others => '0');
                            rs2_internal <=                                  (others => '0');
                            imm_internal <=                                  i_instruction(31 downto 12)                       
                                                                           & "000000000000";
                            
                            -- i_instruction identification
                            case i_instruction(6 downto 2) is

                                when "01101" =>
                                    opcode <= i_LUI; 
                                    illegal_internal2 <= '0';
                                when "00101" =>
                                    opcode <= i_AUIPC; 
                                    illegal_internal2 <= '0';
                                when others =>
                                    opcode <= i_NOP; 
                                    illegal_internal2 <= '1';
                            
                            end case;

                        -- Jumps
                        when J =>
                            rd_internal <=                                  (others => '0');
                            rs1_internal <=                                 i_instruction(19 downto 15); 
                            rs2_internal <=                                 i_instruction(24 downto 20);
                            imm_internal <=                                 (others => i_instruction(31));
                            imm_internal(20 downto 1) <=                    i_instruction(31)                                 
                                                                          & i_instruction(19 downto 12)     
                                                                          & i_instruction(20)                   
                                                                          & i_instruction(30 downto 21);
                            imm_internal(0) <=                              '0';
                            
                            -- i_instruction identification
                            case i_instruction(6 downto 2) is

                                when "11011" =>
                                    opcode <= i_JAL; 
                                    illegal_internal2 <= '0';
                                when others =>
                                    opcode <= i_NOP; 
                                    illegal_internal2 <= '1';
                            
                            end case;

                        when NOP =>
                            rd_internal <=                                  (others => '0');
                            rs1_internal <=                                 (others => '0');
                            rs2_internal <=                                 (others => '0');
                            imm_internal <=                                 (others => '0');
                            opcode <=                                       i_NOP;  
                            illegal_internal2 <=                            '0';                     
                        
                        when others =>
                            rd_internal <=                                  (others => '0');
                            rs1_internal <=                                 (others => '0');
                            rs2_internal <=                                 (others => '0');
                            imm_internal <=                                 (others => '0');
                            opcode <=                                       i_NOP;
                            illegal_internal2 <=                            '1'; 

                    end case;
            
                end if;

            end process;

        -- Compute the illegal status
        illegal_internal_out <= illegal_internal or illegal_internal2;

        -- Output signals, while encouting for illegal state.
        illegal <= illegal_internal_out;

        rs1 <= rs1_internal when illegal_internal_out = '0' else
            std_logic_vector(to_unsigned(0, rs1'length));
        rs2 <= rs2_internal when illegal_internal_out = '0' else
            std_logic_vector(to_unsigned(0, rs2'length));
        rd <= rd_internal when illegal_internal_out = '0' else
            std_logic_vector(to_unsigned(0, rd'length));
        imm <= imm_internal when illegal_internal_out = '0' else
            std_logic_vector(to_unsigned(0, imm'length));

    end architecture;