library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity alu is 
end entity;

architecture behavioral of alu is
    begin
    end architecture;