library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity b_decoder is 
end entity;

architecture behavioral of b_decoder is
    begin
    end architecture;