LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;

ENTITY timer_peripheral_tb IS
END ENTITY;

ARCHITECTURE behavioral OF timer_peripheral_tb IS
BEGIN
END ARCHITECTURE;