LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;

ENTITY serial_peripheral IS
END ENTITY;

ARCHITECTURE behavioral OF serial_peripheral IS
BEGIN
END ARCHITECTURE;