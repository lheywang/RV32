/*
 *  File :      rtl/core/core.sv
 *
 *  Author :    l.heywang <leonard.heywang@proton.me>
 *  Date :      25/10.2025
 *  
 *  Brief :     This file assemble all of the core components into
 *              a single entity, easier to use rather than a lot
 *              of smallers modules.
 */

`timescale 1ns / 1ps

module core (

);

endmodule
