library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity decoder is 
end entity;

architecture behavioral of decoder is
    begin
    end architecture;