LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;

ENTITY ulpi_peripheral IS
END ENTITY;

ARCHITECTURE behavioral OF ulpi_peripheral IS
BEGIN
END ARCHITECTURE;