/*
 *  File :      rtl/core/issuer.sv
 *
 *  Author :    l.heywang <leonard.heywang@proton.me>
 *  Date :      25/10.2025
 *  
 *  Brief :     This file define the issuer module, the one charged to 
 *              split incomming instructions into the right ALU, and start
 *              as many instruction as it can to get the maximal performance
 *              available from the core.
 */

module issuer ();

endmodule
