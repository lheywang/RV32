library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity core_controller_tb is 
end entity;

architecture behavioral of core_controller_tb is
    begin
    end architecture;