library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity pwm_peripheral is 
end entity;

architecture behavioral of pwm_peripheral is
    begin
    end architecture;