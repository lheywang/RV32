--! @file rv32.vhd
--! @brief This is the top entity of the RV32 core, which include peripherals and memories. Theses may be vendor dependant.
--! @author l.heywang <leonard.heywang@proton.me>
--! date 05-10-25

LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;

ENTITY rv32 IS
END ENTITY;

ARCHITECTURE behavioral OF rv32 IS
BEGIN
END ARCHITECTURE;