library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity sdram_tb is 
end entity;

architecture behavioral of sdram_tb is
    begin
    end architecture;