library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity cache is 
end entity;

architecture behavioral of cache is
    begin
    end architecture;