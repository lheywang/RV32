/*
 *  File :      rtl/core/assembly/assembly_alu.sv
 *
 *  Author :    l.heywang <leonard.heywang@proton.me>
 *  Date :      25/10.2025
 *  
 *  Brief :     This file assemble all of the ALU with the issuer
 *              and commiter units. This is done to make the global
 *              core.sv file much more readable.
 */

module assembly_alu (

);

endmodule
