library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity u_decoder is 
end entity;

architecture behavioral of u_decoder is
    begin
    end architecture;