library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity memory is 
end entity;

architecture behavioral of memory is
    begin
    end architecture;