library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity s_decoder is 
end entity;

architecture behavioral of s_decoder is
    begin
    end architecture;