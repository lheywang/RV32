library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity argb_peripheral is 
end entity;

architecture behavioral of argb_peripheral is
    begin
    end architecture;