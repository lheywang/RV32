library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity timer_peripheral_tb is 
end entity;

architecture behavioral of timer_peripheral_tb is
    begin
    end architecture;